// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by rejaz on Sun 31 Jul 18:00:08 PKT 2022
//
// cmd:    swerv -iccm_size=4 -dccm_size=4 -snapshot=4kbmemories 
//

`include "common_defines.vh"
`undef RV_ASSERT_ON
`undef TEC_RV_ICG
`define RV_PHYSICAL 1
